module mongo
