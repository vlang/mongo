module mongo

