module bson

// http://mongoc.org/libbson/current/bson_t.html
pub struct C.bson_t {}

// http://mongoc.org/libbson/current/bson_oid_t.html
pub struct C.bson_oid_t {}

// http://mongoc.org/libbson/current/bson_subtype_t.html
pub struct C.bson_subtype_t {}

// http://mongoc.org/libbson/current/bson_context_t.html
pub struct C.bson_context_t {}

// http://mongoc.org/libbson/current/bson_subtype_t.html
pub struct C.bson_subtyper_t {}

// http://mongoc.org/libbson/current/bson_decimal128_t.html
pub struct C.bson_decimal128_t {}

// http://mongoc.org/libbson/current/bson_iter_t.html
pub struct C.bson_iter_t {}

// http://mongoc.org/libbson/current/bson_value_t.html
pub struct C.bson_value_t {}

// http://mongoc.org/libbson/current/bson_error_t.html
pub struct C.bson_error_t {}