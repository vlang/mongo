module bson

/*
pub fn (value string) bson_type() voidptr
{
	return C.BCON_UTF8(value.str)
}

pub fn (value int) bson_type() voidptr
{
	return C.BSON_APPEND_INT32(value)
}

pub fn (value byte) bson_type() voidptr
{
	return C.BCON_BOOL(value.str)
}

pub fn (value bool) bson_type() voidptr
{
	return C.BCON_BOOL(value.str)
}

pub fn (value Oid) bson_type() voidptr
{
	return C.BCON_OID(values)
}
*/
