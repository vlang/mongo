module mongo

// http://mongoc.org/libmongoc/current/mongoc_client_t.html
pub struct C.mongoc_client_t {}

// http://mongoc.org/libmongoc/current/mongoc_client_pool_new.html
pub struct C.mongoc_client_pool_t {}

// http://mongoc.org/libmongoc/current/mongoc_database_t.html
pub struct C.mongoc_database_t {}

// http://mongoc.org/libmongoc/current/mongoc_collection_t.html
pub struct C.mongoc_collection_t {}

// http://mongoc.org/libmongoc/current/mongoc_write_concern_t.html
pub struct C.mongoc_write_concern_t {}

// http://mongoc.org/libmongoc/current/mongoc_uri_t.html
pub struct C.mongoc_uri_t {}

// http://mongoc.org/libmongoc/current/mongoc_cursor_t.html
pub struct C.mongoc_cursor_t {}

// http://mongoc.org/libmongoc/1.17.0/mongoc_query_flags_t.html
pub struct C.mongoc_query_flags_t {}

// http://mongoc.org/libmongoc/current/mongoc_read_prefs_t.html
pub struct C.mongoc_read_prefs_t {}

// http://mongoc.org/libmongoc/current/mongoc_stream_t.html
pub struct C.mongoc_stream_t {}

// http://mongoc.org/libmongoc/current/mongoc_stream_file_t.html
pub struct C.mongoc_stream_file_t {}
